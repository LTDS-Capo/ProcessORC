module StackCache #(
    parameter 
)(
    input clk,
    input clk_en,
    input sync_rst,

    input                          InstructionValid,
    input                          InstructionIsARunahead, // Potentially already allocated to the Push Queue

    input                          CacheLineInREQ,
    output                         CacheLineInACK,
    input  [CACHELINEBITWIDTH-1:0] CacheLineInData,

    output                         CacheLineOutREQ,
    input                          CacheLineOutACK,
    output [CACHELINEBITWIDTH-1:0] CacheLineOutData,

    input                   [31:0] StackUpperBound,
    input                   [31:0] StackLowerBound,
    input                          StackDirection, // 0 - Grows Down with Push, 1 - Grows Up with Push

    input                   [31:0] StackPointerIn,
    output                  [31:0] StackPointerOut,
    input                          StackPointerSwap, // Force Cache Flush and Fetch


);


    // Push Queue/Wait Table with 4bit Write Tags
    // 16 entry table with a 4 bit tag
    // Tag is generated by a counter that is allowed to wrap around,
    // If Current tag points to a currently in-flight Tag, Stall until condition clears

        //! Have a mechanism to pre-write Pushes to Cache lines that are still being fetched

    // Cache Lines are 8 elements
    // 4 Cache Lines In size

    // 32 entry table to show status of each stack element

// ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~

    // States
        // Normal Operation
        // Prefetch Push - Pre-write to Cache line (Can not happen on speculation)
        // Prefetch Pop
        // Cache Miss on Push - Pre-write to Cache line (Can not happen on speculation)
        // Cache Miss on Pop
        // Cache Flush - Post Swap
        // Cache Fill - Post Swap
    //

    // Stack Pointer
        // Pointer

        // Shadow Pointer

        wire CacheSwap = StackPointerSwap;
    //

    // Speculative Write History

    //

    // Push Wait Table
        StackCache_PushWaitTable_Dynamic #(
            .DATABITWIDTH(DATABITWIDTH)
        ) DynamicWaitTable (
            .clk                         (),
            .clk_en                      (),
            .sync_rst                    (),
            .Speculating                 (),
            .MispredictedSpeculationPulse(),
            .AllowedToSpeculate          (),
            .NoPendingWrites             (),
            .InstructionValid            (),
            .WillBeWriting               (),
            .TagValid                    (),
            .AssignedTag                 (),
            .StackPointer                (),
            .StackWriteEn                (),
            .StackWriteTag               (),
            .WriteAddress                ()
        );
    //

    // Cache Line Generation

    //

    // Stack Cache Entry Status Buffer
        // 4x Vectors, 
    //

endmodule : StackCache

