module BranchTargetBuffer #(
    parameter DATABITWIDTH = 16
)(
    input clk,
    input clk_en,
    input sync_rst,

    input [DATABITWIDTH-1:0] 
);



endmodule : BranchTargetBuffer