module PlatformIndependant_TopLevel (
    ports
);
    


    // Initialization
    // Notes:
    // In:
    // Out:
    
    //

    CPU_TopLevel CPU (

    );
    

    // IO
    // Notes:
    // In:
    // Out:
    
    //


endmodule