module System_TopLevel (
    //ports
);
    
    // Initialization
    // Notes:
    // In:
    // Out:
    
    //

    CPU_TopLevel CPU (

    );
    
endmodule