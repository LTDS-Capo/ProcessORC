Hi! I am AFK for a min, making some tea :)
