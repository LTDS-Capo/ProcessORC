module IOManager #(
    parameter TOTALIOBYTES = 128,
// $PARAMETERS$
    parameter TOTALIOPORTS = 8,
// $ENDPARAMETERS$
)(
    ports
);


// $GEN$ CaseGen([8:Addr, 4:Output], CaseConfig.txt)
// $GENEND$



endmodule